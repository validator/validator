<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML 1.0 Strict//EN"
    "http://www.w3.org/TR/xhtml1/DTD/xhtml1-strict.dtd">
<html xmlns="http://www.w3.org/1999/xhtml" xml:lang="sv" lang="sv">
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8" />
  <title>Dokumentation avseende W3C:s CSS-validerare</title>
  <link rev="made" href="mailto:www-validator-css@w3.org" />
  <link rev="start" href="./" title="Hemsida" />
  <style type="text/css" media="all">
    @import "style/base.css";    
    @import "style/docs.css";    
  </style>
  <meta name="revision" content="$Id$" />
  <!-- SSI Template Version: $Id$ -->
</head>

<body>
  <div id="banner">
   <h1 id="title"><a href="https://www.w3.org/"><img alt="W3C" id="logo" src="https://www.w3.org/assets/logos/w3c-2025/svg/margins/w3c-letters-bg-white.svg" /></a>
   <a href="./"><span>CSS valideringstjänst</span></a></h1>
   <p id="tagline">
     Granska formatmallar ("<span xml:lang="en" lang="en">Check Cascading Style Sheets</span>, CSS) och (X)HTML-dokument med formatmallar
   </p>
  </div>


<div id="main">
<!-- This DIV encapsulates everything in this page - necessary for the positioning -->

<div class="doc">
<h2>Dokumentation om CSS-valideraren</h2>

<p id="skip"></p>

<h3 id="use">Resurser för användare</h3>

<dl>
  <dt><a href="./manual.html">Användarmanual</a></dt>
  <dd>Dokumentation om hur CSS-valideraren kan användas</dd>
  <dt><a href="about.html">Om denna tjänst</a></dt>
  <dd>Information om CSS-valideraren, och svar på allmänna frågor</dd>
  <dt><a href="http://www.websitedev.de/css/validator-faq">
      Vanliga frågor och svar om CSS-validerare (FAQ)
      </a></dt>
  <dd>Svar på vanligt förekommande tekniska frågor.</dd>
</dl>

<h3 id="devel">Resurser för utvecklare</h3>


<dl>
  <dt><a href="DOWNLOAD.html">Ladda ned/installera</a></dt>
  <dd>Hur man hämtar källkoden för CSS-valideraren och kör den,
      antingen från kommandoraden eller som en webb-servlet.</dd>
      
  <dt><a href="README">Utvecklarens README</a></dt>
  <dd>En översikt över programkoden i CSS-valideraren</dd>
      
  <dt><a href="./api.html">Web Service API</a></dt>
  <dd>Dokumentation av SOAP 1.2-gränssnitt mot valideraren</dd>
      
  <dt><a href="https://github.com/w3c/css-validator/issues">Buggar</a> &amp; <a href="https://www.w3.org/Bugs/Public/buglist.cgi?bug_status=__open__;product=CSSValidator">Buggar</a></dt>
  <dd>Kända problem i aktuell version av valideraren, och ett
      gränssnitt med vilket man kan meddela nya buggar och problem.
      Se även <a href="Email.html">anvisningar för hur synpunkter delges</a>.</dd>
</dl>



</div>
</div>
<!-- End of "main" DIV. -->

<ul class="navbar"  id="menu">
  <li><strong><a href="./" title="Hemsida för W3C:s CSS valideringstjänst">Hemsida</a></strong> <span class="hideme">|</span></li>
  <li><a href="about.html" title="Om denna tjänst">Om</a> <span class="hideme">|</span></li>
  <li><a href="DOWNLOAD.html" title="Ladda ned CSS-valideraren">Ladda ned</a> <span class="hideme">|</span></li>
  <li><a href="Email.html" title="Hur man ger synpunkter på denna tjänst">Synpunkter</a> <span class="hideme">|</span></li>
  <li><a href="thanks.html" title="Tack och erkännanden">Tack</a><span class="hideme">|</span></li>
</ul>

<ul id="lang_choice">
     
     <li><a href="documentation.html.bg"
    lang="bg"
    xml:lang="bg"
    hreflang="bg"
    rel="alternate">Български</a></li>
  <li><a href="documentation.html.de"
         lang="de"
         xml:lang="de"
         hreflang="de"
         rel="alternate">Deutsch</a>
     </li>
     
     <li><a href="documentation.html.en"
         lang="en"
         xml:lang="en"
         hreflang="en"
         rel="alternate">English</a>
     </li>
     
     <li><a href="documentation.html.es"
         lang="es"
         xml:lang="es"
         hreflang="es"
         rel="alternate">Español</a>
     </li>
     
     <li><a href="documentation.html.fr"
         lang="fr"
         xml:lang="fr"
         hreflang="fr"
         rel="alternate">Français</a>
     </li>
     
     <li><a href="documentation.html.ko"
         lang="ko"
         xml:lang="ko"
         hreflang="ko"
         rel="alternate">한국어</a>
     </li>
     
     <li><a href="documentation.html.it"
         lang="it"
         xml:lang="it"
         hreflang="it"
         rel="alternate">Italiano</a>
     </li>
     
     <li><a href="documentation.html.nl"
         lang="nl"
         xml:lang="nl"
         hreflang="nl"
         rel="alternate">Nederlands</a>
     </li>
     
     <li><a href="documentation.html.ja"
         lang="ja"
         xml:lang="ja"
         hreflang="ja"
         rel="alternate">日本語</a>
     </li>
     
     <li><a href="documentation.html.pl-PL"
         lang="pl-PL"
         xml:lang="pl-PL"
         hreflang="pl-PL"
         rel="alternate">Polski</a>
     </li>
     
     <li><a href="documentation.html.pt-BR"
         lang="pt-BR"
         xml:lang="pt-BR"
         hreflang="pt-BR"
         rel="alternate">Português</a>
     </li>
     
     <li><a href="documentation.html.ru"
         lang="ru"
         xml:lang="ru"
         hreflang="ru"
         rel="alternate">Русский</a>
     </li>
     
     <li><a href="documentation.html.sv"
         lang="sv"
         xml:lang="sv"
         hreflang="sv"
         rel="alternate">Svenska</a>
     </li>
     
     <li><a href="documentation.html.zh-cn"
         lang="zh-cn"
         xml:lang="zh-cn"
         hreflang="zh-cn"
         rel="alternate">简体中文</a>
     </li>
</ul>



<div id="footer">
<p id="activity_logos">

<a href="https://www.w3.org/Style/CSS/learning" title="Mer information om formatmallar"><img src="images/woolly-icon" alt="CSS" /></a>
</p>

<p id="support_logo">
<a href="https://www.w3.org/donate/">
<img src="https://www.w3.org/QA/Tools/I_heart_validator" alt="I heart Validator logo" title=" Validators Donation Program" />
</a>
</p>

<p class="copyright"><span lang="en" dir="ltr">Copyright &copy; 2025 <a href="https://www.w3.org/">World Wide Web Consortium</a>.<br> <abbr title="World Wide Web Consortium">W3C</abbr><sup>&reg;</sup> <a href="https://www.w3.org/policies/#disclaimers">liability</a>, <a href="https://www.w3.org/policies/#trademarks">trademark</a> and <a rel="license" href="https://www.w3.org/copyright/document-license/" title="W3C Document License">permissive license</a> rules apply.</span></p>

</div>
</body>
</html>


